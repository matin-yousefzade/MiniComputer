module MC_TB_BasicCode2();
  reg [31:0]ClientMemWrite,ClientMemAddr,ClientInsAddr;
  reg [4:0]ClientRegAddr;
  reg [1:0]CWDM,CRDM,CRIM;
  reg Start,InitPC,InitLNO,Clk,Rst;
  reg del,tilde,ccb,pipe,ocb,z,y,x,w,v,u,t,s,r,q,p,o,n,m,l,k,j,i,h,g,f,e,d,c,b,a,backtick,undelrine,hat,csb,backslash,osb,Z,Y,X,W,V,U,T,S,R,Q,P,O,N,M,L,K,J,I,H,G,F,E,D,C,B,A,atsign,question,gt,equal,lt,semicolon,colon,n9,n8,n7,n6,n5,n4,n3,n2,n1,n0,slash,dot,minus,comma,plus,asterisk,cp,op,singlequote,ampersand,percent,dollar,sharp,doublequote,exclamation,space,us,rs,gs,fs,esc,sub,em,can,etb,syn,nak,dc4,dc3,dc2,dc1,dle,si,so,cr,ff,vt,lf,ht,bs,bel,ack,enq,eot,etx,stx,soh,null;
  wire [31:0]ClientMemRead,ClientInsRead,ClientRegRead,WID;
  wire [7:0]CIMRD,AIMRD,Opcode;
  wire [5:0]ps;
  wire [4:0]CPUps;
  wire [3:0]Cps;
  wire Ready,CReady,CPUReady;
  MiniComputer G1(ClientMemWrite,ClientMemAddr,ClientInsAddr,ClientRegAddr,CWDM,CRDM,CRIM,Start,InitPC,InitLNO,Clk,Rst,del,tilde,ccb,pipe,ocb,z,y,x,w,v,u,t,s,r,q,p,o,n,m,l,k,j,i,h,g,f,e,d,c,b,a,backtick,undelrine,hat,csb,backslash,osb,Z,Y,X,W,V,U,T,S,R,Q,P,O,N,M,L,K,J,I,H,G,F,E,D,C,B,A,atsign,question,gt,equal,lt,semicolon,colon,n9,n8,n7,n6,n5,n4,n3,n2,n1,n0,slash,dot,minus,comma,plus,asterisk,cp,op,singlequote,ampersand,percent,dollar,sharp,doublequote,exclamation,space,us,rs,gs,fs,esc,sub,em,can,etb,syn,nak,dc4,dc3,dc2,dc1,dle,si,so,cr,ff,vt,lf,ht,bs,bel,ack,enq,eot,etx,stx,soh,null,ClientMemRead,ClientInsRead,ClientRegRead,WID,CIMRD,AIMRD,Opcode,ps,CPUps,Cps,Ready,CReady,CPUReady);
  initial begin
    Clk=0;
    forever begin
      #50 Clk=!Clk;
    end
  end
  initial begin
    {del,tilde,ccb,pipe,ocb,z,y,x,w,v,u,t,s,r,q,p,o,n,m,l,k,j,i,h,g,f,e,d,c,b,a,backtick,undelrine,hat,csb,backslash,osb,Z,Y,X,W,V,U,T,S,R,Q,P,O,N,M,L,K,J,I,H,G,F,E,D,C,B,A,atsign,question,gt,equal,lt,semicolon,colon,n9,n8,n7,n6,n5,n4,n3,n2,n1,n0,slash,dot,minus,comma,plus,asterisk,cp,op,singlequote,ampersand,percent,dollar,sharp,doublequote,exclamation,space,us,rs,gs,fs,esc,sub,em,can,etb,syn,nak,dc4,dc3,dc2,dc1,dle,si,so,cr,ff,vt,lf,ht,bs,bel,ack,enq,eot,etx,stx,soh,null}=128'h0;
    Start=0;
    Rst=1;
    #100
    Rst=0;
    InitPC=1;
    InitLNO=1;
    #100
    InitPC=0;
    InitLNO=0;
    Start=1;
    #100
    Start=0;
    #100
    //**********************************
    //**********************************
    //**********************************
    //label div
    //label sr
    //num x 8
    //assign R1 I4
    //assign R2 I4
    //beq R1 R2 Lsr
    //div:div R4 I9 R2
    //exit
    //sr:xor R3 Vx R1
    //ror Vx R3 I5
    //jmp Ldiv
    //**********************************
    //**********************************
    //**********************************
    //label div
    l=1;
    #100
    l=0;
    a=1;
    #100
    a=0;
    b=1;
    #100
    b=0;
    e=1;
    #100
    e=0;
    l=1;
    #100
    l=0;
    space=1;
    #100
    space=0;
    d=1;
    #100
    d=0;
    i=1;
    #100
    i=0;
    v=1;
    #100
    v=0;
    lf=1;
    #100
    lf=0;
    //label sr
    l=1;
    #100
    l=0;
    a=1;
    #100
    a=0;
    b=1;
    #100
    b=0;
    e=1;
    #100
    e=0;
    l=1;
    #100
    l=0;
    space=1;
    #100
    space=0;
    s=1;
    #100
    s=0;
    r=1;
    #100
    r=0;
    lf=1;
    #100
    lf=0;
    //num x 8
    n=1;
    #100
    n=0;
    u=1;
    #100
    u=0;
    m=1;
    #100
    m=0;
    space=1;
    #100
    space=0;
    x=1;
    #100
    x=0;
    space=1;
    #100
    space=0;
    n8=1;
    #100
    n8=0;
    lf=1;
    #100
    lf=0;
    //assign R1 I4
    a=1;
    #100
    a=0;
    s=1;
    #100
    #100
    s=0;
    i=1;
    #100
    i=0;
    g=1;
    #100
    g=0;
    n=1;
    #100
    n=0;
    space=1;
    #100
    space=0;
    R=1;
    #100
    R=0;
    n1=1;
    #100
    n1=0;
    space=1;
    #100
    space=0;
    I=1;
    #100
    I=0;
    n4=1;
    #100
    n4=0;
    lf=1;
    #100
    lf=0;
    //assign R2 I4
    a=1;
    #100
    a=0;
    s=1;
    #100
    #100
    s=0;
    i=1;
    #100
    i=0;
    g=1;
    #100
    g=0;
    n=1;
    #100
    n=0;
    space=1;
    #100
    space=0;
    R=1;
    #100
    R=0;
    n2=1;
    #100
    n2=0;
    space=1;
    #100
    space=0;
    I=1;
    #100
    I=0;
    n4=1;
    #100
    n4=0;
    lf=1;
    #100
    lf=0;
    //beq R1 R2 Lsr
    b=1;
    #100
    b=0;
    e=1;
    #100
    e=0;
    q=1;
    #100
    q=0;
    space=1;
    #100
    space=0;
    R=1;
    #100
    R=0;
    n1=1;
    #100
    n1=0;
    space=1;
    #100
    space=0;
    R=1;
    #100
    R=0;
    n2=1;
    #100
    n2=0;
    space=1;
    #100
    space=0;
    L=1;
    #100
    L=0;
    s=1;
    #100
    s=0;
    r=1;
    #100
    r=0;
    lf=1;
    #100
    lf=0;
    //div:div R4 I9 R2
    d=1;
    #100
    d=0;
    i=1;
    #100
    i=0;
    v=1;
    #100
    v=0;
    colon=1;
    #100
    colon=0;
    d=1;
    #100
    d=0;
    i=1;
    #100
    i=0;
    v=1;
    #100
    v=0;
    space=1;
    #100
    space=0;
    R=1;
    #100
    R=0;
    n4=1;
    #100
    n4=0;
    space=1;
    #100
    space=0;
    I=1;
    #100
    I=0;
    n9=1;
    #100
    n9=0;
    space=1;
    #100
    space=0;
    R=1;
    #100
    R=0;
    n2=1;
    #100
    n2=0;
    lf=1;
    #100
    lf=0;
    //exit
    e=1;
    #100
    e=0;
    x=1;
    #100
    x=0;
    i=1;
    #100
    i=0;
    t=1;
    #100
    t=0;
    lf=1;
    #100
    lf=0;
    //sr:xor R3 Vx R1
    s=1;
    #100
    s=0;
    r=1;
    #100
    r=0;
    colon=1;
    #100
    colon=0;
    x=1;
    #100
    x=0;
    o=1;
    #100
    o=0;
    r=1;
    #100
    r=0;
    space=1;
    #100
    space=0;
    R=1;
    #100
    R=0;
    n3=1;
    #100
    n3=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    x=1;
    #100
    x=0;
    space=1;
    #100
    space=0;
    R=1;
    #100
    R=0;
    n1=1;
    #100
    n1=0;
    lf=1;
    #100
    lf=0;
    //ror Vx R3 I5
    r=1;
    #100
    r=0;
    o=1;
    #100
    o=0;
    r=1;
    #100
    r=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    x=1;
    #100
    x=0;
    space=1;
    #100
    space=0;
    R=1;
    #100
    R=0;
    n3=1;
    #100
    n3=0;
    space=1;
    #100
    space=0;
    I=1;
    #100
    I=0;
    n5=1;
    #100
    n5=0;
    lf=1;
    #100
    lf=0;
    //jmp Ldiv
    j=1;
    #100
    j=0;
    m=1;
    #100
    m=0;
    p=1;
    #100
    p=0;
    space=1;
    #100
    space=0;
    L=1;
    #100
    L=0;
    d=1;
    #100
    d=0;
    i=1;
    #100
    i=0;
    v=1;
    #100
    v=0;
    etx=1;
    #10000000
    ClientInsAddr=32'h0;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h4;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h8;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'hC;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h10;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h14;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h18;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h1C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h20;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h24;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h28;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h2C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h30;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h34;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h38;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h3C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h40;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h44;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h48;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h4C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h50;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h54;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h58;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h5C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h60;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h64;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h68;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h6C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h70;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h74;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h78;
    CRIM=2'h3;
    #107
    ClientInsAddr=32'h7C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h80;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h84;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h88;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h8C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h90;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h94;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h98;
    CRIM=2'h3;
    #107
    ClientInsAddr=32'h9C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'hA0;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'hA4;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'hA8;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'hAC;
    CRIM=2'h3;
    #100
    CRIM=2'h0;
    //************************************
    //************************************
    //************************************
    ClientRegAddr=5'h1;
    #100
    ClientRegAddr=5'h2;
    #100
    ClientRegAddr=5'h3;
    #100
    ClientRegAddr=5'h4;
    #100
    //************************************
    //************************************
    //************************************
    ClientMemAddr=32'h8000;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8001;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8002;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8003;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8004;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8005;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8006;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8007;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8008;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8009;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800A;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800B;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800C;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800D;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800E;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800F;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8010;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8011;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8012;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8013;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8014;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8015;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8016;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8017;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8018;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8019;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801A;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801B;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801C;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801D;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801E;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801F;
    CRDM=2'h1;
    #100
    $stop;
  end
endmodule