module MiniComputer(input [31:0]ClientMemWrite,ClientMemAddr,ClientInsAddr,input [4:0]ClientRegAddr,input [1:0]CWDM,CRDM,CRIM,input Start,InitPC,InitLNO,Clk,Rst,input del,tilde,ccb,pipe,ocb,z,y,x,w,v,u,t,s,r,q,p,o,n,m,l,k,j,i,h,g,f,e,d,c,b,a,backtick,undelrine,hat,csb,backslash,osb,Z,Y,X,W,V,U,T,S,R,Q,P,O,N,M,L,K,J,I,H,G,F,E,D,C,B,A,atsign,question,gt,equal,lt,semicolon,colon,n9,n8,n7,n6,n5,n4,n3,n2,n1,n0,slash,dot,minus,comma,plus,asterisk,cp,op,singlequote,ampersand,percent,dollar,sharp,doublequote,exclamation,space,us,rs,gs,fs,esc,sub,em,can,etb,syn,nak,dc4,dc3,dc2,dc1,dle,si,so,cr,ff,vt,lf,ht,bs,bel,ack,enq,eot,etx,stx,soh,null,output [31:0]ClientMemRead,ClientInsRead,ClientRegRead,WID,output [7:0]CIMRD,AIMRD,Opcode,output [5:0]ps,output [4:0]CPUps,output [3:0]Cps,output Ready,CReady,CPUReady);
  wire [127:0]other;
  wire [31:0]MemWriteBus,MemAddrBus,MemReadBus,WIA;
  wire [15:0]CIMA,CIMR;
  wire [8:0]AIMA;
  wire [7:0]CIMWD;
  wire [4:0]AIMUnity;
  wire [3:0]ParIPP,IPP;
  wire [2:0]grt;
  wire [1:0]WIM,WDMB,RDMB,ParTR;
  wire ETXF,InitETXF,LdETXF,XF,InitXF,LdXF,ParIFR,LdIFR,LdTR,InitCIMR,LdCIMR,CIPP,InitIPP,ParLdIPP,CCIM,InitCIM,ParLdCIM,CAIM;
  wire InitAIM,PAK,WCIM,RCIM,WAIM,RAIM,Co1,Co2,Co3,CStart,OCStart,VCStart,CPUStart,AStart,VMgrt,IOACgrt,VCgrt,CPUgrt,OCReady,VCReady,VCHalfReady;
  wire VMreq,IOACreq,VCreq,CPUreq,CLNO,InitAIM2;
  Register_1b_Init R1(1'h1,Clk,Rst,InitETXF,LdETXF,ETXF);
  Register_1b_Init R2(1'h1,Clk,Rst,InitXF,LdXF,XF);
  Register_16b_Init R3(CIMA,Clk,Rst,InitCIMR,LdCIMR,CIMR);
  Counter_4b_Par C1(ParIPP,CIPP,InitIPP,ParLdIPP,Clk,Rst,IPP,Co1);
  Counter_5b C2(CAIM,InitAIM,Clk,Rst,AIMUnity,Co2);
  Counter_16b_Par C3(CIMR,CCIM,InitCIM,ParLdCIM,Clk,Rst,CIMA,Co3);
  Adder_9b G1({IPP,5'h0},{4'h0,AIMUnity},AIMA);
  Keyboard G2(other,del,tilde,ccb,pipe,ocb,z,y,x,w,v,u,t,s,r,q,p,o,n,m,l,k,j,i,h,g,f,e,d,c,b,a,backtick,undelrine,hat,csb,backslash,osb,Z,Y,X,W,V,U,T,S,R,Q,P,O,N,M,L,K,J,I,H,G,F,E,D,C,B,A,atsign,question,gt,equal,lt,semicolon,colon,n9,n8,n7,n6,n5,n4,n3,n2,n1,n0,slash,dot,minus,comma,plus,asterisk,cp,op,singlequote,ampersand,percent,dollar,sharp,doublequote,exclamation,space,us,rs,gs,fs,esc,sub,em,can,etb,syn,nak,dc4,dc3,dc2,dc1,dle,si,so,cr,ff,vt,lf,ht,bs,bel,ack,enq,eot,etx,stx,soh,null,CIMWD,PAK);
  ClientInstructionMemory G3(CIMA,CIMWD,WCIM,RCIM,Clk,Rst,CIMRD);
  AloneInstructionMemory G4(AIMA,CIMRD,WAIM,RAIM,InitAIM2,Clk,Rst,AIMRD);
  DataMemory G5(MemWriteBus,MemAddrBus,ClientMemWrite,ClientMemAddr,WDMB,RDMB,CWDM,CRDM,Clk,Rst,MemReadBus,ClientMemRead);
  Compiler G6(WIA,MemReadBus,AIMRD,Opcode,IPP,CStart,VMgrt,IOACgrt,Clk,Rst,WID,MemWriteBus,MemAddrBus,Cps,WDMB,RDMB,WIM,CReady,VMreq,IOACreq,CLNO);
  VariableCreator G7(MemReadBus,AIMRD,ParTR,VCStart,ParIFR,LdTR,LdIFR,VCgrt,Clk,Rst,MemWriteBus,MemAddrBus,WDMB,RDMB,VCReady,VCHalfReady,VCreq);
  CPU G8(WID,ClientInsRead,ClientInsAddr,MemReadBus,ClientRegAddr,WIM,CRIM,CPUStart,InitPC,InitLNO,CLNO,CPUgrt,Clk,Rst,ClientRegRead,WIA,MemWriteBus,MemAddrBus,CPUps,WDMB,RDMB,CPUReady,CPUreq);
  OpcodeConvertor G9(AIMRD,OCStart,Clk,Rst,Opcode,OCReady);
  Arbiter G10({3'h0,VMreq,IOACreq,VCreq,CPUreq},AStart,Clk,Rst,{grt,VMgrt,IOACgrt,VCgrt,CPUgrt});
  MC_Controller G11(Opcode,CIMWD,CIMRD,AIMRD,IPP,Start,PAK,ETXF,XF,CReady,OCReady,VCHalfReady,VCReady,CPUReady,Clk,Rst,ps,ParIPP,ParTR,Ready,InitCIMR,LdCIMR,InitETXF,LdETXF,InitXF,LdXF,ParIFR,LdIFR,LdTR,WCIM,RCIM,CCIM,InitCIM,ParLdCIM,WAIM,RAIM,CAIM,InitAIM,CIPP,InitIPP,ParLdIPP,CStart,OCStart,VCStart,CPUStart,AStart,InitAIM2);
endmodule



module MC_TB_PrimeNumber();
  reg [31:0]ClientMemWrite,ClientMemAddr,ClientInsAddr;
  reg [4:0]ClientRegAddr;
  reg [1:0]CWDM,CRDM,CRIM;
  reg Start,InitPC,InitLNO,Clk,Rst;
  reg del,tilde,ccb,pipe,ocb,z,y,x,w,v,u,t,s,r,q,p,o,n,m,l,k,j,i,h,g,f,e,d,c,b,a,backtick,undelrine,hat,csb,backslash,osb,Z,Y,X,W,V,U,T,S,R,Q,P,O,N,M,L,K,J,I,H,G,F,E,D,C,B,A,atsign,question,gt,equal,lt,semicolon,colon,n9,n8,n7,n6,n5,n4,n3,n2,n1,n0,slash,dot,minus,comma,plus,asterisk,cp,op,singlequote,ampersand,percent,dollar,sharp,doublequote,exclamation,space,us,rs,gs,fs,esc,sub,em,can,etb,syn,nak,dc4,dc3,dc2,dc1,dle,si,so,cr,ff,vt,lf,ht,bs,bel,ack,enq,eot,etx,stx,soh,null;
  wire [31:0]ClientMemRead,ClientInsRead,ClientRegRead,WID;
  wire [7:0]CIMRD,AIMRD,Opcode;
  wire [5:0]ps;
  wire [4:0]CPUps;
  wire [3:0]Cps;
  wire Ready,CReady,CPUReady;
  MiniComputer G1(ClientMemWrite,ClientMemAddr,ClientInsAddr,ClientRegAddr,CWDM,CRDM,CRIM,Start,InitPC,InitLNO,Clk,Rst,del,tilde,ccb,pipe,ocb,z,y,x,w,v,u,t,s,r,q,p,o,n,m,l,k,j,i,h,g,f,e,d,c,b,a,backtick,undelrine,hat,csb,backslash,osb,Z,Y,X,W,V,U,T,S,R,Q,P,O,N,M,L,K,J,I,H,G,F,E,D,C,B,A,atsign,question,gt,equal,lt,semicolon,colon,n9,n8,n7,n6,n5,n4,n3,n2,n1,n0,slash,dot,minus,comma,plus,asterisk,cp,op,singlequote,ampersand,percent,dollar,sharp,doublequote,exclamation,space,us,rs,gs,fs,esc,sub,em,can,etb,syn,nak,dc4,dc3,dc2,dc1,dle,si,so,cr,ff,vt,lf,ht,bs,bel,ack,enq,eot,etx,stx,soh,null,ClientMemRead,ClientInsRead,ClientRegRead,WID,CIMRD,AIMRD,Opcode,ps,CPUps,Cps,Ready,CReady,CPUReady);
  initial begin
    Clk=0;
    forever begin
      #50 Clk=!Clk;
    end
  end
  initial begin
    {del,tilde,ccb,pipe,ocb,z,y,x,w,v,u,t,s,r,q,p,o,n,m,l,k,j,i,h,g,f,e,d,c,b,a,backtick,undelrine,hat,csb,backslash,osb,Z,Y,X,W,V,U,T,S,R,Q,P,O,N,M,L,K,J,I,H,G,F,E,D,C,B,A,atsign,question,gt,equal,lt,semicolon,colon,n9,n8,n7,n6,n5,n4,n3,n2,n1,n0,slash,dot,minus,comma,plus,asterisk,cp,op,singlequote,ampersand,percent,dollar,sharp,doublequote,exclamation,space,us,rs,gs,fs,esc,sub,em,can,etb,syn,nak,dc4,dc3,dc2,dc1,dle,si,so,cr,ff,vt,lf,ht,bs,bel,ack,enq,eot,etx,stx,soh,null}=128'h0;
    Start=0;
    Rst=1;
    #100
    Rst=0;
    InitPC=1;
    InitLNO=1;
    #100
    InitPC=0;
    InitLNO=0;
    Start=1;
    #100
    Start=0;
    #100
    //**********************************
    //**********************************
    //**********************************
    //label Loop
    //label CNL
    //num x 35
    //num i 2
    //num pn 1
    //num y
    //Loop:div Vy Vx Vi
    //mlt Vy Vy Vi
    //beq Vx Vy LCNL
    //add Vi Vi I1
    //blt Vi Vx LLoop
    //exit
    //CNL:assign Vpn I0
    //exit
    //**********************************
    //**********************************
    //**********************************
    //label Loop
    l=1;
    #100
    l=0;
    a=1;
    #100
    a=0;
    b=1;
    #100
    b=0;
    e=1;
    #100
    e=0;
    l=1;
    #100
    l=0;
    space=1;
    #100
    space=0;
    L=1;
    #100
    L=0;
    o=1;
    #100
    #100
    o=0;
    p=1;
    #100
    p=0;
    lf=1;
    #100
    lf=0;
    //label CNL
    l=1;
    #100
    l=0;
    a=1;
    #100
    a=0;
    b=1;
    #100
    b=0;
    e=1;
    #100
    e=0;
    l=1;
    #100
    l=0;
    space=1;
    #100
    space=0;
    C=1;
    #100
    C=0;
    N=1;
    #100
    N=0;
    L=1;
    #100
    L=0;
    lf=1;
    #100
    lf=0;
    //num x 35
    n=1;
    #100
    n=0;
    u=1;
    #100
    u=0;
    m=1;
    #100
    m=0;
    space=1;
    #100
    space=0;
    x=1;
    #100
    x=0;
    space=1;
    #100
    space=0;
    n3=1;
    #100
    n3=0;
    n5=1;
    #100
    n5=0;
    lf=1;
    #100
    lf=0;
    //num i 2
    n=1;
    #100
    n=0;
    u=1;
    #100
    u=0;
    m=1;
    #100
    m=0;
    space=1;
    #100
    space=0;
    i=1;
    #100
    i=0;
    space=1;
    #100
    space=0;
    n2=1;
    #100
    n2=0;
    lf=1;
    #100
    lf=0;
    //num pn 1
    n=1;
    #100
    n=0;
    u=1;
    #100
    u=0;
    m=1;
    #100
    m=0;
    space=1;
    #100
    space=0;
    p=1;
    #100
    p=0;
    n=1;
    #100
    n=0;
    space=1;
    #100
    space=0;
    n1=1;
    #100
    n1=0;
    lf=1;
    #100
    lf=0;
    //num y
    n=1;
    #100
    n=0;
    u=1;
    #100
    u=0;
    m=1;
    #100
    m=0;
    space=1;
    #100
    space=0;
    y=1;
    #100
    y=0;
    lf=1;
    #100
    lf=0;
    //Loop:div Vy Vx Vi
    L=1;
    #100
    L=0;
    o=1;
    #100
    #100
    o=0;
    p=1;
    #100
    p=0;
    colon=1;
    #100
    colon=0;
    d=1;
    #100
    d=0;
    i=1;
    #100
    i=0;
    v=1;
    #100
    v=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    y=1;
    #100
    y=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    x=1;
    #100
    x=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    i=1;
    #100
    i=0;
    lf=1;
    #100
    lf=0;
    //mlt Vy Vy Vi
    m=1;
    #100
    m=0;
    l=1;
    #100
    l=0;
    t=1;
    #100
    t=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    y=1;
    #100
    y=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    y=1;
    #100
    y=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    i=1;
    #100
    i=0;
    lf=1;
    #100
    lf=0;
    //beq Vx Vy LCNL
    b=1;
    #100
    b=0;
    e=1;
    #100
    e=0;
    q=1;
    #100
    q=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    x=1;
    #100
    x=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    y=1;
    #100
    y=0;
    space=1;
    #100
    space=0;
    L=1;
    #100
    L=0;
    C=1;
    #100
    C=0;
    N=1;
    #100
    N=0;
    L=1;
    #100
    L=0;
    lf=1;
    #100
    lf=0;
    //add Vi Vi I1
    a=1;
    #100
    a=0;
    d=1;
    #100
    #100
    d=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    i=1;
    #100
    i=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    i=1;
    #100
    i=0;
    space=1;
    #100
    space=0;
    I=1;
    #100
    I=0;
    n1=1;
    #100
    n1=0;
    lf=1;
    #100
    lf=0;
    //blt Vi Vx LLoop
    b=1;
    #100
    b=0;
    l=1;
    #100
    l=0;
    t=1;
    #100
    t=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    i=1;
    #100
    i=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    x=1;
    #100
    x=0;
    space=1;
    #100
    space=0;
    L=1;
    #100
    #100
    L=0;
    o=1;
    #100
    #100
    o=0;
    p=1;
    #100
    p=0;
    lf=1;
    #100
    lf=0;
    //exit
    e=1;
    #100
    e=0;
    x=1;
    #100
    x=0;
    i=1;
    #100
    i=0;
    t=1;
    #100
    t=0;
    lf=1;
    #100
    lf=0;
    //CNL:assign Vpn I0
    C=1;
    #100
    C=0;
    N=1;
    #100
    N=0;
    L=1;
    #100
    L=0;
    colon=1;
    #100
    colon=0;
    a=1;
    #100
    a=0;
    s=1;
    #100
    #100
    s=0;
    i=1;
    #100
    i=0;
    g=1;
    #100
    g=0;
    n=1;
    #100
    n=0;
    space=1;
    #100
    space=0;
    V=1;
    #100
    V=0;
    p=1;
    #100
    p=0;
    n=1;
    #100
    n=0;
    space=1;
    #100
    space=0;
    I=1;
    #100
    I=0;
    n0=1;
    #100
    n0=0;
    lf=1;
    #100
    lf=0;
    //exit
    e=1;
    #100
    e=0;
    x=1;
    #100
    x=0;
    i=1;
    #100
    i=0;
    t=1;
    #100
    t=0;
    etx=1;
    #10000000
    ClientInsAddr=32'h0;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h4;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h8;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'hC;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h10;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h14;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h18;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h1C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h20;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h24;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h28;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h2C;
    CRIM=2'h3;
    #100  
    ClientInsAddr=32'h30;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h34;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h38;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h3C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h40;
    CRIM=2'h3;
    #100  
    ClientInsAddr=32'h44;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h48;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h4C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h50;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h54;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h58;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h5C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h60;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h64;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h68;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h6C;
    CRIM=2'h3;
    #100  
    ClientInsAddr=32'h70;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h74;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h78;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h7C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h80;
    CRIM=2'h3;
    #100  
    ClientInsAddr=32'h84;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h88;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h8C;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h90;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h94;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h98;
    CRIM=2'h3;
    #100
    ClientInsAddr=32'h9C;
    CRIM=2'h3;
    #100
    CRIM=2'h0;
    //************************************
    //************************************
    //************************************
    ClientMemAddr=32'h8000;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8001;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8002;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8003;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8004;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8005;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8006;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8007;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8008;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8009;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800A;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800B;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800C;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800D;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800E;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h800F;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8010;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8011;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8012;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8013;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8014;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8015;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8016;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8017;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8018;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8019;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801A;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801B;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801C;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801D;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801E;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h801F;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8020;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8021;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8022;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8023;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8024;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8025;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8026;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8027;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8028;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8029;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h802A;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h802B;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h802C;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h802D;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h802E;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h802F;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8030;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8031;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8032;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8033;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8034;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8035;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8036;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8037;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8038;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h8039;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h803A;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h803B;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h803C;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h803D;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h803E;
    CRDM=2'h1;
    #100
    ClientMemAddr=32'h803F;
    CRDM=2'h1;
    #100
    $stop;
  end
endmodule