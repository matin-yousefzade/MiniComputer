module Plus4(input [31:0]A,output [31:0]W);
  assign W=A+4;
endmodule