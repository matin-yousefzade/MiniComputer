module Subtractor_3b(input [2:0]A,B,output [2:0]W);
  assign W=A-B;
endmodule