module Inc_3b(input [2:0]A,output [2:0]W);
  assign W=A+1;
endmodule


module Inc_2b(input [1:0]A,output [1:0]W);
  assign W=A+1;
endmodule